--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
-- All globally shared constants are defined in this package.                       +
--                                                                                  +
-- File : glbSharedTypes.vhd                                                        +
--+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;
use IEEE.math_real.all;

package glbSharedTypes is

	constant   FU_ADDRESS_W    : integer   := 6;
	constant   FU_DATA_W       : integer   := 5;
	constant   FU_FIFO_IDX_W   : integer   := 1; 
	constant   FU_INPUT_W      : integer   := (2 ** FU_DATA_W)-1;
	
	-- Memory element constants. If there are multiple memory elements, first $MEM_SELECT_BITLENGTH bits
	-- of $MEM_ADDR_LENGTH are used for memory unit selection.
	-- Every unit has $BANK_SIZE long,word addressable flat address space.
	-- At this stage, number of load and store units are the same.
	constant   MEM_WORD_LENGTH	   	: integer   := 32;	--Number of bytes in each word
	constant   MEM_NR_ELEMENTS	   	: integer   := 4;		--Number of load and store elements(for each)
	constant   MEM_BANK_SIZE	   	: integer   := 64;	--Memory size in 4-byte words
	constant   MEM_ADDR_LENGTH   		: integer   := integer(log2(REAL(MEM_NR_ELEMENTS * MEM_BANK_SIZE)));
	constant   MEM_SELECT_BITLENGTH 	: integer 	:= integer(log2(REAL(MEM_NR_ELEMENTS)));
	
	type ram_type is array (0 to MEM_BANK_SIZE - 1) of std_logic_vector (MEM_WORD_LENGTH - 1 downto 0);
	
	type sorterIOVector_t is record
		--vld		: std_logic;												-- Validity assertion register bits
		tarAddr	: std_logic_vector(FU_ADDRESS_W  -1 downto 0);	-- target FU address ( The validity of address is encapsulated in the msb of the tarAddr (Active Low) VALD=0, INVD=1 )
		srcAddr	: std_logic_vector(FU_ADDRESS_W  -2 downto 0);	-- source FU address 
		data	: std_logic_vector(FU_DATA_W     -1 downto 0);	-- data to be routed
		fifoIdx	: std_logic_vector(FU_FIFO_IDX_W -1 downto 0);	-- Input fifo index
	end record;
	
	type validVector_t is array ( 0 to FU_INPUT_W ) of std_logic;

	-- IO wires for the network
	type bitonStageBus_t is array (0 to FU_INPUT_W) of sorterIOVector_t;
	-- Invalid address table
	type invAddArr_t is array ( 0 to FU_INPUT_W) of std_logic_vector (FU_ADDRESS_W-2 downto 0);
	-- DTN-Routing table type
	type dtnRoutTbl_t is array (0 to FU_INPUT_W,0 to FU_INPUT_W) of std_logic_vector(FU_ADDRESS_W  -2 downto 0);
	-- DTN-Router states
	type dtnRouterStates_t is (DETERMINE ,ROUTE, LOCKED ) ;
	
	constant InvAddr : invAddArr_t := (	"00000","00001","00010","00011","00100","00101","00110","00111",
													"01000","01001","01010","01011","01100","01101","01110","01111",
													"10000","10001","10010","10011","10100","10101","10110","10111",
													"11000","11001","11010","11011","11100","11101","11110","11111");
	-- Reset values for pipeline stage registers												
	constant pRegDefVal	: bitonStageBus_t := ( others => ("000000","00000", "00000","0"));
	-- Reset values for DTN-Router ports
	constant dtnRtrDefVal: sorterIOVector_t := ("000000","00000", "00000","0");
	-- Forward routing table
	constant FW_RT: dtnRoutTbl_t:=(("00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111"),
											("00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ),
											("00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ),
											("00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ),
											("00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ),
											("00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ),
											("00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ),
											("00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ),
											("01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ),
											("01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ),
											("01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ),
											("01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ),
											("01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ),
											("01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ),
											("01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ),
											("01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ),
											("10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ),
											("10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ),
											("10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ),
											("10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ),
											("10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ),
											("10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ),
											("10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ),
											("10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ),
											("11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ),
											("11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ),
											("11010" ,"11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ),
											("11011" ,"11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ),
											("11100" ,"11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ),
											("11101" ,"11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ),
											("11110" ,"11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ),
											("11111" ,"00000" ,"00001" ,"00010" ,"00011" ,"00100" ,"00101" ,"00110" ,"00111" ,"01000" ,"01001" ,"01010" ,"01011" ,"01100" ,"01101" ,"01110" ,"01111" ,"10000" ,"10001" ,"10010" ,"10011" ,"10100" ,"10101" ,"10110" ,"10111" ,"11000" ,"11001" ,"11010" ,"11011" ,"11100" ,"11101" ,"11110" ));
	-- Reverse routing table
	constant RV_RT: dtnRoutTbl_t:=(("11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000"),
											("11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ),
											("11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ),
											("11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ),
											("11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ),
											("11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ),
											("11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ),
											("11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ),
											("10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ),
											("10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ),
											("10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ),
											("10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ),
											("10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ),
											("10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ),
											("10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ),
											("10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ),
											("01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ),
											("01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ),
											("01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ),
											("01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ),
											("01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ),
											("01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ),
											("01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ),
											("01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ),
											("00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ),
											("00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ),
											("00101" ,"00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ),
											("00100" ,"00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ),
											("00011" ,"00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ),
											("00010" ,"00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ),
											("00001" ,"00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ),
											("00000" ,"11111" ,"11110" ,"11101" ,"11100" ,"11011" ,"11010" ,"11001" ,"11000" ,"10111" ,"10110" ,"10101" ,"10100" ,"10011" ,"10010" ,"10001" ,"10000" ,"01111" ,"01110" ,"01101" ,"01100" ,"01011" ,"01010" ,"01001" ,"01000" ,"00111" ,"00110" ,"00101" ,"00100" ,"00011" ,"00010" ,"00001" ));

	-- fucntion reuturns the validity the given address
	function isAddrValid(addr : IN std_logic_vector (FU_ADDRESS_W  -1 downto 0)) return std_logic;
	function getAddressIdx(addr : IN std_logic_vector (FU_ADDRESS_W  -1 downto 0)) return integer;
end glbSharedTypes;



package body glbSharedTypes is
	-- returns true if the address is VALID else returns false
	function isAddrValid(addr : IN std_logic_vector (FU_ADDRESS_W  -1 downto 0)) return std_logic is
	begin
		return not (addr(FU_ADDRESS_W  -1));
	end function isAddrValid;

	function getAddressIdx(addr : IN std_logic_vector (FU_ADDRESS_W  -1 downto 0)) return integer is
	begin
		return to_integer(unsigned(addr));
	end function getAddressIdx;	
	
end glbSharedTypes;
